/*************************************************
* Copyright 2024 NTT Corporation, FUJITSU LIMITED
* Licensed under the Apache License, Version 2.0, see LICENSE for details.
* SPDX-License-Identifier: Apache-2.0
*************************************************/

`timescale 1ns/100ps
`default_nettype none

module chain_control (
    input wire ap_clk,
    input wire ap_rst_n,
    output wire detect_fault,
    output wire interrupt,
    output wire [63:0] m_axi_extif0_buffer_rd_ARADDR,
    output wire [1:0] m_axi_extif0_buffer_rd_ARBURST,
    output wire [3:0] m_axi_extif0_buffer_rd_ARCACHE,
    output wire [0:0] m_axi_extif0_buffer_rd_ARID,
    output wire [7:0] m_axi_extif0_buffer_rd_ARLEN,
    output wire [1:0] m_axi_extif0_buffer_rd_ARLOCK,
    output wire [2:0] m_axi_extif0_buffer_rd_ARPROT,
    output wire [3:0] m_axi_extif0_buffer_rd_ARQOS,
    input wire m_axi_extif0_buffer_rd_ARREADY,
    output wire [3:0] m_axi_extif0_buffer_rd_ARREGION,
    output wire [2:0] m_axi_extif0_buffer_rd_ARSIZE,
    output wire m_axi_extif0_buffer_rd_ARVALID,
    output wire [63:0] m_axi_extif0_buffer_rd_AWADDR,
    output wire [1:0] m_axi_extif0_buffer_rd_AWBURST,
    output wire [3:0] m_axi_extif0_buffer_rd_AWCACHE,
    output wire [0:0] m_axi_extif0_buffer_rd_AWID,
    output wire [7:0] m_axi_extif0_buffer_rd_AWLEN,
    output wire [1:0] m_axi_extif0_buffer_rd_AWLOCK,
    output wire [2:0] m_axi_extif0_buffer_rd_AWPROT,
    output wire [3:0] m_axi_extif0_buffer_rd_AWQOS,
    input wire m_axi_extif0_buffer_rd_AWREADY,
    output wire [3:0] m_axi_extif0_buffer_rd_AWREGION,
    output wire [2:0] m_axi_extif0_buffer_rd_AWSIZE,
    output wire m_axi_extif0_buffer_rd_AWVALID,
    input wire [0:0] m_axi_extif0_buffer_rd_BID,
    output wire m_axi_extif0_buffer_rd_BREADY,
    input wire [1:0] m_axi_extif0_buffer_rd_BRESP,
    input wire m_axi_extif0_buffer_rd_BVALID,
    input wire [511:0] m_axi_extif0_buffer_rd_RDATA,
    input wire [0:0] m_axi_extif0_buffer_rd_RID,
    input wire m_axi_extif0_buffer_rd_RLAST,
    output wire m_axi_extif0_buffer_rd_RREADY,
    input wire [1:0] m_axi_extif0_buffer_rd_RRESP,
    input wire m_axi_extif0_buffer_rd_RVALID,
    output wire [511:0] m_axi_extif0_buffer_rd_WDATA,
    output wire [0:0] m_axi_extif0_buffer_rd_WID,
    output wire m_axi_extif0_buffer_rd_WLAST,
    input wire m_axi_extif0_buffer_rd_WREADY,
    output wire [63:0] m_axi_extif0_buffer_rd_WSTRB,
    output wire m_axi_extif0_buffer_rd_WVALID,
    output wire [63:0] m_axi_extif0_buffer_wr_ARADDR,
    output wire [1:0] m_axi_extif0_buffer_wr_ARBURST,
    output wire [3:0] m_axi_extif0_buffer_wr_ARCACHE,
    output wire [0:0] m_axi_extif0_buffer_wr_ARID,
    output wire [7:0] m_axi_extif0_buffer_wr_ARLEN,
    output wire [1:0] m_axi_extif0_buffer_wr_ARLOCK,
    output wire [2:0] m_axi_extif0_buffer_wr_ARPROT,
    output wire [3:0] m_axi_extif0_buffer_wr_ARQOS,
    input wire m_axi_extif0_buffer_wr_ARREADY,
    output wire [3:0] m_axi_extif0_buffer_wr_ARREGION,
    output wire [2:0] m_axi_extif0_buffer_wr_ARSIZE,
    output wire m_axi_extif0_buffer_wr_ARVALID,
    output wire [63:0] m_axi_extif0_buffer_wr_AWADDR,
    output wire [1:0] m_axi_extif0_buffer_wr_AWBURST,
    output wire [3:0] m_axi_extif0_buffer_wr_AWCACHE,
    output wire [0:0] m_axi_extif0_buffer_wr_AWID,
    output wire [7:0] m_axi_extif0_buffer_wr_AWLEN,
    output wire [1:0] m_axi_extif0_buffer_wr_AWLOCK,
    output wire [2:0] m_axi_extif0_buffer_wr_AWPROT,
    output wire [3:0] m_axi_extif0_buffer_wr_AWQOS,
    input wire m_axi_extif0_buffer_wr_AWREADY,
    output wire [3:0] m_axi_extif0_buffer_wr_AWREGION,
    output wire [2:0] m_axi_extif0_buffer_wr_AWSIZE,
    output wire m_axi_extif0_buffer_wr_AWVALID,
    input wire [0:0] m_axi_extif0_buffer_wr_BID,
    output wire m_axi_extif0_buffer_wr_BREADY,
    input wire [1:0] m_axi_extif0_buffer_wr_BRESP,
    input wire m_axi_extif0_buffer_wr_BVALID,
    input wire [511:0] m_axi_extif0_buffer_wr_RDATA,
    input wire [0:0] m_axi_extif0_buffer_wr_RID,
    input wire m_axi_extif0_buffer_wr_RLAST,
    output wire m_axi_extif0_buffer_wr_RREADY,
    input wire [1:0] m_axi_extif0_buffer_wr_RRESP,
    input wire m_axi_extif0_buffer_wr_RVALID,
    output wire [511:0] m_axi_extif0_buffer_wr_WDATA,
    output wire [0:0] m_axi_extif0_buffer_wr_WID,
    output wire m_axi_extif0_buffer_wr_WLAST,
    input wire m_axi_extif0_buffer_wr_WREADY,
    output wire [63:0] m_axi_extif0_buffer_wr_WSTRB,
    output wire m_axi_extif0_buffer_wr_WVALID,
    output wire [63:0] m_axi_extif1_buffer_rd_ARADDR,
    output wire [1:0] m_axi_extif1_buffer_rd_ARBURST,
    output wire [3:0] m_axi_extif1_buffer_rd_ARCACHE,
    output wire [0:0] m_axi_extif1_buffer_rd_ARID,
    output wire [7:0] m_axi_extif1_buffer_rd_ARLEN,
    output wire [1:0] m_axi_extif1_buffer_rd_ARLOCK,
    output wire [2:0] m_axi_extif1_buffer_rd_ARPROT,
    output wire [3:0] m_axi_extif1_buffer_rd_ARQOS,
    input wire m_axi_extif1_buffer_rd_ARREADY,
    output wire [3:0] m_axi_extif1_buffer_rd_ARREGION,
    output wire [2:0] m_axi_extif1_buffer_rd_ARSIZE,
    output wire m_axi_extif1_buffer_rd_ARVALID,
    output wire [63:0] m_axi_extif1_buffer_rd_AWADDR,
    output wire [1:0] m_axi_extif1_buffer_rd_AWBURST,
    output wire [3:0] m_axi_extif1_buffer_rd_AWCACHE,
    output wire [0:0] m_axi_extif1_buffer_rd_AWID,
    output wire [7:0] m_axi_extif1_buffer_rd_AWLEN,
    output wire [1:0] m_axi_extif1_buffer_rd_AWLOCK,
    output wire [2:0] m_axi_extif1_buffer_rd_AWPROT,
    output wire [3:0] m_axi_extif1_buffer_rd_AWQOS,
    input wire m_axi_extif1_buffer_rd_AWREADY,
    output wire [3:0] m_axi_extif1_buffer_rd_AWREGION,
    output wire [2:0] m_axi_extif1_buffer_rd_AWSIZE,
    output wire m_axi_extif1_buffer_rd_AWVALID,
    input wire [0:0] m_axi_extif1_buffer_rd_BID,
    output wire m_axi_extif1_buffer_rd_BREADY,
    input wire [1:0] m_axi_extif1_buffer_rd_BRESP,
    input wire m_axi_extif1_buffer_rd_BVALID,
    input wire [511:0] m_axi_extif1_buffer_rd_RDATA,
    input wire [0:0] m_axi_extif1_buffer_rd_RID,
    input wire m_axi_extif1_buffer_rd_RLAST,
    output wire m_axi_extif1_buffer_rd_RREADY,
    input wire [1:0] m_axi_extif1_buffer_rd_RRESP,
    input wire m_axi_extif1_buffer_rd_RVALID,
    output wire [511:0] m_axi_extif1_buffer_rd_WDATA,
    output wire [0:0] m_axi_extif1_buffer_rd_WID,
    output wire m_axi_extif1_buffer_rd_WLAST,
    input wire m_axi_extif1_buffer_rd_WREADY,
    output wire [63:0] m_axi_extif1_buffer_rd_WSTRB,
    output wire m_axi_extif1_buffer_rd_WVALID,
    output wire [63:0] m_axi_extif1_buffer_wr_ARADDR,
    output wire [1:0] m_axi_extif1_buffer_wr_ARBURST,
    output wire [3:0] m_axi_extif1_buffer_wr_ARCACHE,
    output wire [0:0] m_axi_extif1_buffer_wr_ARID,
    output wire [7:0] m_axi_extif1_buffer_wr_ARLEN,
    output wire [1:0] m_axi_extif1_buffer_wr_ARLOCK,
    output wire [2:0] m_axi_extif1_buffer_wr_ARPROT,
    output wire [3:0] m_axi_extif1_buffer_wr_ARQOS,
    input wire m_axi_extif1_buffer_wr_ARREADY,
    output wire [3:0] m_axi_extif1_buffer_wr_ARREGION,
    output wire [2:0] m_axi_extif1_buffer_wr_ARSIZE,
    output wire m_axi_extif1_buffer_wr_ARVALID,
    output wire [63:0] m_axi_extif1_buffer_wr_AWADDR,
    output wire [1:0] m_axi_extif1_buffer_wr_AWBURST,
    output wire [3:0] m_axi_extif1_buffer_wr_AWCACHE,
    output wire [0:0] m_axi_extif1_buffer_wr_AWID,
    output wire [7:0] m_axi_extif1_buffer_wr_AWLEN,
    output wire [1:0] m_axi_extif1_buffer_wr_AWLOCK,
    output wire [2:0] m_axi_extif1_buffer_wr_AWPROT,
    output wire [3:0] m_axi_extif1_buffer_wr_AWQOS,
    input wire m_axi_extif1_buffer_wr_AWREADY,
    output wire [3:0] m_axi_extif1_buffer_wr_AWREGION,
    output wire [2:0] m_axi_extif1_buffer_wr_AWSIZE,
    output wire m_axi_extif1_buffer_wr_AWVALID,
    input wire [0:0] m_axi_extif1_buffer_wr_BID,
    output wire m_axi_extif1_buffer_wr_BREADY,
    input wire [1:0] m_axi_extif1_buffer_wr_BRESP,
    input wire m_axi_extif1_buffer_wr_BVALID,
    input wire [511:0] m_axi_extif1_buffer_wr_RDATA,
    input wire [0:0] m_axi_extif1_buffer_wr_RID,
    input wire m_axi_extif1_buffer_wr_RLAST,
    output wire m_axi_extif1_buffer_wr_RREADY,
    input wire [1:0] m_axi_extif1_buffer_wr_RRESP,
    input wire m_axi_extif1_buffer_wr_RVALID,
    output wire [511:0] m_axi_extif1_buffer_wr_WDATA,
    output wire [0:0] m_axi_extif1_buffer_wr_WID,
    output wire m_axi_extif1_buffer_wr_WLAST,
    input wire m_axi_extif1_buffer_wr_WREADY,
    output wire [63:0] m_axi_extif1_buffer_wr_WSTRB,
    output wire m_axi_extif1_buffer_wr_WVALID,
    output wire [63:0] m_axis_egr_rx_resp_TDATA,
    input wire m_axis_egr_rx_resp_TREADY,
    output wire m_axis_egr_rx_resp_TVALID,
    output wire [63:0] m_axis_extif0_cmd_TDATA,
    input wire m_axis_extif0_cmd_TREADY,
    output wire m_axis_extif0_cmd_TVALID,
    output wire [63:0] m_axis_extif1_cmd_TDATA,
    input wire m_axis_extif1_cmd_TREADY,
    output wire m_axis_extif1_cmd_TVALID,
    output wire [511:0] m_axis_ingr_tx_data_TDATA,
    input wire m_axis_ingr_tx_data_TREADY,
    output wire m_axis_ingr_tx_data_TVALID,
    output wire [63:0] m_axis_ingr_tx_req_TDATA,
    input wire m_axis_ingr_tx_req_TREADY,
    output wire m_axis_ingr_tx_req_TVALID,
    input wire [11:0] s_axi_control_ARADDR,
    output wire s_axi_control_ARREADY,
    input wire s_axi_control_ARVALID,
    input wire [11:0] s_axi_control_AWADDR,
    output wire s_axi_control_AWREADY,
    input wire s_axi_control_AWVALID,
    input wire s_axi_control_BREADY,
    output wire [1:0] s_axi_control_BRESP,
    output wire s_axi_control_BVALID,
    output wire [31:0] s_axi_control_RDATA,
    input wire s_axi_control_RREADY,
    output wire [1:0] s_axi_control_RRESP,
    output wire s_axi_control_RVALID,
    input wire [31:0] s_axi_control_WDATA,
    output wire s_axi_control_WREADY,
    input wire [3:0] s_axi_control_WSTRB,
    input wire s_axi_control_WVALID,
    input wire [511:0] s_axis_egr_rx_data_TDATA,
    output wire s_axis_egr_rx_data_TREADY,
    input wire s_axis_egr_rx_data_TVALID,
    input wire [63:0] s_axis_egr_rx_req_TDATA,
    output wire s_axis_egr_rx_req_TREADY,
    input wire s_axis_egr_rx_req_TVALID,
    input wire [127:0] s_axis_extif0_evt_TDATA,
    output wire s_axis_extif0_evt_TREADY,
    input wire s_axis_extif0_evt_TVALID,
    input wire [127:0] s_axis_extif1_evt_TDATA,
    output wire s_axis_extif1_evt_TREADY,
    input wire s_axis_extif1_evt_TVALID,
    input wire [63:0] s_axis_ingr_tx_resp_TDATA,
    output wire s_axis_ingr_tx_resp_TREADY,
    input wire s_axis_ingr_tx_resp_TVALID
);

  assign interrupt = 1'b0;
  
  wire[9:0] w_streamif_stall;
  assign w_streamif_stall[0] = m_axis_ingr_tx_req_TVALID  & ~ m_axis_ingr_tx_req_TREADY;
  assign w_streamif_stall[1] = s_axis_ingr_tx_resp_TVALID & ~ s_axis_ingr_tx_resp_TREADY;
  assign w_streamif_stall[2] = m_axis_ingr_tx_data_TVALID & ~ m_axis_ingr_tx_data_TREADY;
  assign w_streamif_stall[3] = s_axis_egr_rx_req_TVALID   & ~ s_axis_egr_rx_req_TREADY;
  assign w_streamif_stall[4] = m_axis_egr_rx_resp_TVALID  & ~ m_axis_egr_rx_resp_TREADY;
  assign w_streamif_stall[5] = s_axis_egr_rx_data_TVALID  & ~ s_axis_egr_rx_data_TREADY;
  assign w_streamif_stall[6] = s_axis_extif0_evt_TVALID   & ~ s_axis_extif0_evt_TREADY;
  assign w_streamif_stall[7] = m_axis_extif0_cmd_TVALID   & ~ m_axis_extif0_cmd_TREADY;
  assign w_streamif_stall[8] = s_axis_extif1_evt_TVALID   & ~ s_axis_extif1_evt_TREADY;
  assign w_streamif_stall[9] = m_axis_extif1_cmd_TVALID   & ~ m_axis_extif1_cmd_TREADY;

  chain_control_bd chain_control_bd_i (
      .ap_clk(ap_clk),
      .ap_rst_n(ap_rst_n),
      .detect_fault(detect_fault),
      .m_axi_extif0_buffer_rd_araddr(m_axi_extif0_buffer_rd_ARADDR),
      .m_axi_extif0_buffer_rd_arburst(m_axi_extif0_buffer_rd_ARBURST),
      .m_axi_extif0_buffer_rd_arcache(m_axi_extif0_buffer_rd_ARCACHE),
      .m_axi_extif0_buffer_rd_arid(m_axi_extif0_buffer_rd_ARID),
      .m_axi_extif0_buffer_rd_arlen(m_axi_extif0_buffer_rd_ARLEN),
      .m_axi_extif0_buffer_rd_arlock(m_axi_extif0_buffer_rd_ARLOCK),
      .m_axi_extif0_buffer_rd_arprot(m_axi_extif0_buffer_rd_ARPROT),
      .m_axi_extif0_buffer_rd_arqos(m_axi_extif0_buffer_rd_ARQOS),
      .m_axi_extif0_buffer_rd_arready(m_axi_extif0_buffer_rd_ARREADY),
      .m_axi_extif0_buffer_rd_arregion(m_axi_extif0_buffer_rd_ARREGION),
      .m_axi_extif0_buffer_rd_arsize(m_axi_extif0_buffer_rd_ARSIZE),
      .m_axi_extif0_buffer_rd_arvalid(m_axi_extif0_buffer_rd_ARVALID),
      .m_axi_extif0_buffer_rd_awaddr(m_axi_extif0_buffer_rd_AWADDR),
      .m_axi_extif0_buffer_rd_awburst(m_axi_extif0_buffer_rd_AWBURST),
      .m_axi_extif0_buffer_rd_awcache(m_axi_extif0_buffer_rd_AWCACHE),
      .m_axi_extif0_buffer_rd_awid(m_axi_extif0_buffer_rd_AWID),
      .m_axi_extif0_buffer_rd_awlen(m_axi_extif0_buffer_rd_AWLEN),
      .m_axi_extif0_buffer_rd_awlock(m_axi_extif0_buffer_rd_AWLOCK),
      .m_axi_extif0_buffer_rd_awprot(m_axi_extif0_buffer_rd_AWPROT),
      .m_axi_extif0_buffer_rd_awqos(m_axi_extif0_buffer_rd_AWQOS),
      .m_axi_extif0_buffer_rd_awready(m_axi_extif0_buffer_rd_AWREADY),
      .m_axi_extif0_buffer_rd_awregion(m_axi_extif0_buffer_rd_AWREGION),
      .m_axi_extif0_buffer_rd_awsize(m_axi_extif0_buffer_rd_AWSIZE),
      .m_axi_extif0_buffer_rd_awvalid(m_axi_extif0_buffer_rd_AWVALID),
      .m_axi_extif0_buffer_rd_bid(m_axi_extif0_buffer_rd_BID),
      .m_axi_extif0_buffer_rd_bready(m_axi_extif0_buffer_rd_BREADY),
      .m_axi_extif0_buffer_rd_bresp(m_axi_extif0_buffer_rd_BRESP),
      .m_axi_extif0_buffer_rd_bvalid(m_axi_extif0_buffer_rd_BVALID),
      .m_axi_extif0_buffer_rd_rdata(m_axi_extif0_buffer_rd_RDATA),
      .m_axi_extif0_buffer_rd_rid(m_axi_extif0_buffer_rd_RID),
      .m_axi_extif0_buffer_rd_rlast(m_axi_extif0_buffer_rd_RLAST),
      .m_axi_extif0_buffer_rd_rready(m_axi_extif0_buffer_rd_RREADY),
      .m_axi_extif0_buffer_rd_rresp(m_axi_extif0_buffer_rd_RRESP),
      .m_axi_extif0_buffer_rd_rvalid(m_axi_extif0_buffer_rd_RVALID),
      .m_axi_extif0_buffer_rd_wdata(m_axi_extif0_buffer_rd_WDATA),
      .m_axi_extif0_buffer_rd_wid(m_axi_extif0_buffer_rd_WID),
      .m_axi_extif0_buffer_rd_wlast(m_axi_extif0_buffer_rd_WLAST),
      .m_axi_extif0_buffer_rd_wready(m_axi_extif0_buffer_rd_WREADY),
      .m_axi_extif0_buffer_rd_wstrb(m_axi_extif0_buffer_rd_WSTRB),
      .m_axi_extif0_buffer_rd_wvalid(m_axi_extif0_buffer_rd_WVALID),
      .m_axi_extif0_buffer_wr_araddr(m_axi_extif0_buffer_wr_ARADDR),
      .m_axi_extif0_buffer_wr_arburst(m_axi_extif0_buffer_wr_ARBURST),
      .m_axi_extif0_buffer_wr_arcache(m_axi_extif0_buffer_wr_ARCACHE),
      .m_axi_extif0_buffer_wr_arid(m_axi_extif0_buffer_wr_ARID),
      .m_axi_extif0_buffer_wr_arlen(m_axi_extif0_buffer_wr_ARLEN),
      .m_axi_extif0_buffer_wr_arlock(m_axi_extif0_buffer_wr_ARLOCK),
      .m_axi_extif0_buffer_wr_arprot(m_axi_extif0_buffer_wr_ARPROT),
      .m_axi_extif0_buffer_wr_arqos(m_axi_extif0_buffer_wr_ARQOS),
      .m_axi_extif0_buffer_wr_arready(m_axi_extif0_buffer_wr_ARREADY),
      .m_axi_extif0_buffer_wr_arregion(m_axi_extif0_buffer_wr_ARREGION),
      .m_axi_extif0_buffer_wr_arsize(m_axi_extif0_buffer_wr_ARSIZE),
      .m_axi_extif0_buffer_wr_arvalid(m_axi_extif0_buffer_wr_ARVALID),
      .m_axi_extif0_buffer_wr_awaddr(m_axi_extif0_buffer_wr_AWADDR),
      .m_axi_extif0_buffer_wr_awburst(m_axi_extif0_buffer_wr_AWBURST),
      .m_axi_extif0_buffer_wr_awcache(m_axi_extif0_buffer_wr_AWCACHE),
      .m_axi_extif0_buffer_wr_awid(m_axi_extif0_buffer_wr_AWID),
      .m_axi_extif0_buffer_wr_awlen(m_axi_extif0_buffer_wr_AWLEN),
      .m_axi_extif0_buffer_wr_awlock(m_axi_extif0_buffer_wr_AWLOCK),
      .m_axi_extif0_buffer_wr_awprot(m_axi_extif0_buffer_wr_AWPROT),
      .m_axi_extif0_buffer_wr_awqos(m_axi_extif0_buffer_wr_AWQOS),
      .m_axi_extif0_buffer_wr_awready(m_axi_extif0_buffer_wr_AWREADY),
      .m_axi_extif0_buffer_wr_awregion(m_axi_extif0_buffer_wr_AWREGION),
      .m_axi_extif0_buffer_wr_awsize(m_axi_extif0_buffer_wr_AWSIZE),
      .m_axi_extif0_buffer_wr_awvalid(m_axi_extif0_buffer_wr_AWVALID),
      .m_axi_extif0_buffer_wr_bid(m_axi_extif0_buffer_wr_BID),
      .m_axi_extif0_buffer_wr_bready(m_axi_extif0_buffer_wr_BREADY),
      .m_axi_extif0_buffer_wr_bresp(m_axi_extif0_buffer_wr_BRESP),
      .m_axi_extif0_buffer_wr_bvalid(m_axi_extif0_buffer_wr_BVALID),
      .m_axi_extif0_buffer_wr_rdata(m_axi_extif0_buffer_wr_RDATA),
      .m_axi_extif0_buffer_wr_rid(m_axi_extif0_buffer_wr_RID),
      .m_axi_extif0_buffer_wr_rlast(m_axi_extif0_buffer_wr_RLAST),
      .m_axi_extif0_buffer_wr_rready(m_axi_extif0_buffer_wr_RREADY),
      .m_axi_extif0_buffer_wr_rresp(m_axi_extif0_buffer_wr_RRESP),
      .m_axi_extif0_buffer_wr_rvalid(m_axi_extif0_buffer_wr_RVALID),
      .m_axi_extif0_buffer_wr_wdata(m_axi_extif0_buffer_wr_WDATA),
      .m_axi_extif0_buffer_wr_wid(m_axi_extif0_buffer_wr_WID),
      .m_axi_extif0_buffer_wr_wlast(m_axi_extif0_buffer_wr_WLAST),
      .m_axi_extif0_buffer_wr_wready(m_axi_extif0_buffer_wr_WREADY),
      .m_axi_extif0_buffer_wr_wstrb(m_axi_extif0_buffer_wr_WSTRB),
      .m_axi_extif0_buffer_wr_wvalid(m_axi_extif0_buffer_wr_WVALID),
      .m_axi_extif1_buffer_rd_araddr(m_axi_extif1_buffer_rd_ARADDR),
      .m_axi_extif1_buffer_rd_arburst(m_axi_extif1_buffer_rd_ARBURST),
      .m_axi_extif1_buffer_rd_arcache(m_axi_extif1_buffer_rd_ARCACHE),
      .m_axi_extif1_buffer_rd_arid(m_axi_extif1_buffer_rd_ARID),
      .m_axi_extif1_buffer_rd_arlen(m_axi_extif1_buffer_rd_ARLEN),
      .m_axi_extif1_buffer_rd_arlock(m_axi_extif1_buffer_rd_ARLOCK),
      .m_axi_extif1_buffer_rd_arprot(m_axi_extif1_buffer_rd_ARPROT),
      .m_axi_extif1_buffer_rd_arqos(m_axi_extif1_buffer_rd_ARQOS),
      .m_axi_extif1_buffer_rd_arready(m_axi_extif1_buffer_rd_ARREADY),
      .m_axi_extif1_buffer_rd_arregion(m_axi_extif1_buffer_rd_ARREGION),
      .m_axi_extif1_buffer_rd_arsize(m_axi_extif1_buffer_rd_ARSIZE),
      .m_axi_extif1_buffer_rd_arvalid(m_axi_extif1_buffer_rd_ARVALID),
      .m_axi_extif1_buffer_rd_awaddr(m_axi_extif1_buffer_rd_AWADDR),
      .m_axi_extif1_buffer_rd_awburst(m_axi_extif1_buffer_rd_AWBURST),
      .m_axi_extif1_buffer_rd_awcache(m_axi_extif1_buffer_rd_AWCACHE),
      .m_axi_extif1_buffer_rd_awid(m_axi_extif1_buffer_rd_AWID),
      .m_axi_extif1_buffer_rd_awlen(m_axi_extif1_buffer_rd_AWLEN),
      .m_axi_extif1_buffer_rd_awlock(m_axi_extif1_buffer_rd_AWLOCK),
      .m_axi_extif1_buffer_rd_awprot(m_axi_extif1_buffer_rd_AWPROT),
      .m_axi_extif1_buffer_rd_awqos(m_axi_extif1_buffer_rd_AWQOS),
      .m_axi_extif1_buffer_rd_awready(m_axi_extif1_buffer_rd_AWREADY),
      .m_axi_extif1_buffer_rd_awregion(m_axi_extif1_buffer_rd_AWREGION),
      .m_axi_extif1_buffer_rd_awsize(m_axi_extif1_buffer_rd_AWSIZE),
      .m_axi_extif1_buffer_rd_awvalid(m_axi_extif1_buffer_rd_AWVALID),
      .m_axi_extif1_buffer_rd_bid(m_axi_extif1_buffer_rd_BID),
      .m_axi_extif1_buffer_rd_bready(m_axi_extif1_buffer_rd_BREADY),
      .m_axi_extif1_buffer_rd_bresp(m_axi_extif1_buffer_rd_BRESP),
      .m_axi_extif1_buffer_rd_bvalid(m_axi_extif1_buffer_rd_BVALID),
      .m_axi_extif1_buffer_rd_rdata(m_axi_extif1_buffer_rd_RDATA),
      .m_axi_extif1_buffer_rd_rid(m_axi_extif1_buffer_rd_RID),
      .m_axi_extif1_buffer_rd_rlast(m_axi_extif1_buffer_rd_RLAST),
      .m_axi_extif1_buffer_rd_rready(m_axi_extif1_buffer_rd_RREADY),
      .m_axi_extif1_buffer_rd_rresp(m_axi_extif1_buffer_rd_RRESP),
      .m_axi_extif1_buffer_rd_rvalid(m_axi_extif1_buffer_rd_RVALID),
      .m_axi_extif1_buffer_rd_wdata(m_axi_extif1_buffer_rd_WDATA),
      .m_axi_extif1_buffer_rd_wid(m_axi_extif1_buffer_rd_WID),
      .m_axi_extif1_buffer_rd_wlast(m_axi_extif1_buffer_rd_WLAST),
      .m_axi_extif1_buffer_rd_wready(m_axi_extif1_buffer_rd_WREADY),
      .m_axi_extif1_buffer_rd_wstrb(m_axi_extif1_buffer_rd_WSTRB),
      .m_axi_extif1_buffer_rd_wvalid(m_axi_extif1_buffer_rd_WVALID),
      .m_axi_extif1_buffer_wr_araddr(m_axi_extif1_buffer_wr_ARADDR),
      .m_axi_extif1_buffer_wr_arburst(m_axi_extif1_buffer_wr_ARBURST),
      .m_axi_extif1_buffer_wr_arcache(m_axi_extif1_buffer_wr_ARCACHE),
      .m_axi_extif1_buffer_wr_arid(m_axi_extif1_buffer_wr_ARID),
      .m_axi_extif1_buffer_wr_arlen(m_axi_extif1_buffer_wr_ARLEN),
      .m_axi_extif1_buffer_wr_arlock(m_axi_extif1_buffer_wr_ARLOCK),
      .m_axi_extif1_buffer_wr_arprot(m_axi_extif1_buffer_wr_ARPROT),
      .m_axi_extif1_buffer_wr_arqos(m_axi_extif1_buffer_wr_ARQOS),
      .m_axi_extif1_buffer_wr_arready(m_axi_extif1_buffer_wr_ARREADY),
      .m_axi_extif1_buffer_wr_arregion(m_axi_extif1_buffer_wr_ARREGION),
      .m_axi_extif1_buffer_wr_arsize(m_axi_extif1_buffer_wr_ARSIZE),
      .m_axi_extif1_buffer_wr_arvalid(m_axi_extif1_buffer_wr_ARVALID),
      .m_axi_extif1_buffer_wr_awaddr(m_axi_extif1_buffer_wr_AWADDR),
      .m_axi_extif1_buffer_wr_awburst(m_axi_extif1_buffer_wr_AWBURST),
      .m_axi_extif1_buffer_wr_awcache(m_axi_extif1_buffer_wr_AWCACHE),
      .m_axi_extif1_buffer_wr_awid(m_axi_extif1_buffer_wr_AWID),
      .m_axi_extif1_buffer_wr_awlen(m_axi_extif1_buffer_wr_AWLEN),
      .m_axi_extif1_buffer_wr_awlock(m_axi_extif1_buffer_wr_AWLOCK),
      .m_axi_extif1_buffer_wr_awprot(m_axi_extif1_buffer_wr_AWPROT),
      .m_axi_extif1_buffer_wr_awqos(m_axi_extif1_buffer_wr_AWQOS),
      .m_axi_extif1_buffer_wr_awready(m_axi_extif1_buffer_wr_AWREADY),
      .m_axi_extif1_buffer_wr_awregion(m_axi_extif1_buffer_wr_AWREGION),
      .m_axi_extif1_buffer_wr_awsize(m_axi_extif1_buffer_wr_AWSIZE),
      .m_axi_extif1_buffer_wr_awvalid(m_axi_extif1_buffer_wr_AWVALID),
      .m_axi_extif1_buffer_wr_bid(m_axi_extif1_buffer_wr_BID),
      .m_axi_extif1_buffer_wr_bready(m_axi_extif1_buffer_wr_BREADY),
      .m_axi_extif1_buffer_wr_bresp(m_axi_extif1_buffer_wr_BRESP),
      .m_axi_extif1_buffer_wr_bvalid(m_axi_extif1_buffer_wr_BVALID),
      .m_axi_extif1_buffer_wr_rdata(m_axi_extif1_buffer_wr_RDATA),
      .m_axi_extif1_buffer_wr_rid(m_axi_extif1_buffer_wr_RID),
      .m_axi_extif1_buffer_wr_rlast(m_axi_extif1_buffer_wr_RLAST),
      .m_axi_extif1_buffer_wr_rready(m_axi_extif1_buffer_wr_RREADY),
      .m_axi_extif1_buffer_wr_rresp(m_axi_extif1_buffer_wr_RRESP),
      .m_axi_extif1_buffer_wr_rvalid(m_axi_extif1_buffer_wr_RVALID),
      .m_axi_extif1_buffer_wr_wdata(m_axi_extif1_buffer_wr_WDATA),
      .m_axi_extif1_buffer_wr_wid(m_axi_extif1_buffer_wr_WID),
      .m_axi_extif1_buffer_wr_wlast(m_axi_extif1_buffer_wr_WLAST),
      .m_axi_extif1_buffer_wr_wready(m_axi_extif1_buffer_wr_WREADY),
      .m_axi_extif1_buffer_wr_wstrb(m_axi_extif1_buffer_wr_WSTRB),
      .m_axi_extif1_buffer_wr_wvalid(m_axi_extif1_buffer_wr_WVALID),
      .m_axis_egr_rx_resp_tdata(m_axis_egr_rx_resp_TDATA),
      .m_axis_egr_rx_resp_tready(m_axis_egr_rx_resp_TREADY),
      .m_axis_egr_rx_resp_tvalid(m_axis_egr_rx_resp_TVALID),
      .m_axis_extif0_cmd_tdata(m_axis_extif0_cmd_TDATA),
      .m_axis_extif0_cmd_tready(m_axis_extif0_cmd_TREADY),
      .m_axis_extif0_cmd_tvalid(m_axis_extif0_cmd_TVALID),
      .m_axis_extif1_cmd_tdata(m_axis_extif1_cmd_TDATA),
      .m_axis_extif1_cmd_tready(m_axis_extif1_cmd_TREADY),
      .m_axis_extif1_cmd_tvalid(m_axis_extif1_cmd_TVALID),
      .m_axis_ingr_tx_data_tdata(m_axis_ingr_tx_data_TDATA),
      .m_axis_ingr_tx_data_tready(m_axis_ingr_tx_data_TREADY),
      .m_axis_ingr_tx_data_tvalid(m_axis_ingr_tx_data_TVALID),
      .m_axis_ingr_tx_req_tdata(m_axis_ingr_tx_req_TDATA),
      .m_axis_ingr_tx_req_tready(m_axis_ingr_tx_req_TREADY),
      .m_axis_ingr_tx_req_tvalid(m_axis_ingr_tx_req_TVALID),
      .s_axi_control_araddr(s_axi_control_ARADDR),
      .s_axi_control_arready(s_axi_control_ARREADY),
      .s_axi_control_arvalid(s_axi_control_ARVALID),
      .s_axi_control_awaddr(s_axi_control_AWADDR),
      .s_axi_control_awready(s_axi_control_AWREADY),
      .s_axi_control_awvalid(s_axi_control_AWVALID),
      .s_axi_control_bready(s_axi_control_BREADY),
      .s_axi_control_bresp(s_axi_control_BRESP),
      .s_axi_control_bvalid(s_axi_control_BVALID),
      .s_axi_control_rdata(s_axi_control_RDATA),
      .s_axi_control_rready(s_axi_control_RREADY),
      .s_axi_control_rresp(s_axi_control_RRESP),
      .s_axi_control_rvalid(s_axi_control_RVALID),
      .s_axi_control_wdata(s_axi_control_WDATA),
      .s_axi_control_wready(s_axi_control_WREADY),
      .s_axi_control_wstrb(s_axi_control_WSTRB),
      .s_axi_control_wvalid(s_axi_control_WVALID),
      .s_axis_egr_rx_data_tdata(s_axis_egr_rx_data_TDATA),
      .s_axis_egr_rx_data_tready(s_axis_egr_rx_data_TREADY),
      .s_axis_egr_rx_data_tvalid(s_axis_egr_rx_data_TVALID),
      .s_axis_egr_rx_req_tdata(s_axis_egr_rx_req_TDATA),
      .s_axis_egr_rx_req_tready(s_axis_egr_rx_req_TREADY),
      .s_axis_egr_rx_req_tvalid(s_axis_egr_rx_req_TVALID),
      .s_axis_extif0_evt_tdata(s_axis_extif0_evt_TDATA),
      .s_axis_extif0_evt_tready(s_axis_extif0_evt_TREADY),
      .s_axis_extif0_evt_tvalid(s_axis_extif0_evt_TVALID),
      .s_axis_extif1_evt_tdata(s_axis_extif1_evt_TDATA),
      .s_axis_extif1_evt_tready(s_axis_extif1_evt_TREADY),
      .s_axis_extif1_evt_tvalid(s_axis_extif1_evt_TVALID),
      .s_axis_ingr_tx_resp_tdata(s_axis_ingr_tx_resp_TDATA),
      .s_axis_ingr_tx_resp_tready(s_axis_ingr_tx_resp_TREADY),
      .s_axis_ingr_tx_resp_tvalid(s_axis_ingr_tx_resp_TVALID),
      .streamif_stall(w_streamif_stall)
  );

endmodule

`default_nettype wire
